Physical Examination||(?:^[\t ]*PHYSICAL EXAMINATION):?[\t \r]*\n
History of Present Illness||(?:^[\t ]*(?:HISTORY OF (?:THE )?(?:PRESENT |PHYSICAL )?ILLNESS)(?: \(HPI(?:, PROBLEM BY PROBLEM)?\))?):?[\t \r]*\n
Past Medical History||(?:^[\t ]*(?:(?:HISTORY OF (?:THE )?PAST ILLNESS)|(?:PAST MEDICAL HISTORY))):?[\t \r]*\n
Chief Complaint||(?:^[\t ]*(?:CHIEF|PRIMARY) COMPLAINTS?):?[\t \r]*\n
Personal and Social History||(?:^[\t ]*(?:(?:PERSONAL (?:(?:AND )?SOCIAL )?HISTORY)?|(?:(?:PSYCHO)?SOC(?:IAL)? HISTORY)|(?:HISTORY (?:OF )(?:OTHER )?SOCIAL (?:FUNCTIONs?|FACTORS?))|(?:PSO)|(?:P?SHX))):?[\t \r]*\n
Review of Systems||(?:^[\t ]*REVIEW OF SYSTEMS?):?[\t \r]*\n
Family Medical History||(?:^[\t ]*(?:FAMILY (?:MEDICAL )?HISTORY)|(?:HISTORY (?:OF )?FAMILY MEMBER DISEASES?)|(?:FAM HX)|FH|FMH|FMHX|FHX):?[\t \r]*\n
Medications||(?:^[\t ]*(?:CURRENT )?MEDICATION)S?:?[\t \r]*\n
Allergies||(?:^[\t ]*ALLERGIES):?[\t \r]*\n
General Exam||(?:^[\t ]*(?:REVIEW (?:OF )?)?GENERAL (?:PHYSICAL )?(?:EXAM(?:INATION)?|STATUS|APPEARANCE|CONSTITUTIONAL)S?(?: SYMPTOMS?)?):?[\t \r]*\n
Vital Signs||(?:^[\t ]*VITAL SIGNS):?[\t \r]*\n
Identifying Data||(?:^[\t ]*IDENTIFYING DATA):?[\t \r]*\n
Clinical History||(?:^[\t ]*CLINICAL HISTORY):?[\t \r]*\n
Current Health||(?:^[\t ]*CURRENT HEALTH(?: STATUS)?):?[\t \r]*\n
Narrative History||(?:^[\t ]*NARRATIVE HISTORY):?[\t \r]*\n
Analysis of Problem||(?:^[\t ]*ANALYSIS (?:OF )?(?:ADMIT(?:TING)? |IDENTIF(?:Y|IED) )?PROBLEMS?):?[\t \r]*\n
Telemetry||(?:^[\t ]*TELE(?:METRY)?):?[\t \r]*\n
Technical Comment||(?:^[\t ]*TECHNICAL COMMENT):?[\t \r]*\n
Discharge Activity||(?:^[\t ]*DISCHARGE ACTIVITY):?[\t \r]*\n
Occupational Environmental History||(?:^[\t ]*OCCUPATION(?:AL)? ENVIRONMENT(?:AL)? HISTORY):?[\t \r]*\n
Immunosuppressants Medications||(?:^[\t ]*(?:CYTOTOXIC )?IMMUNOSUPPRESSANTS? MEDICATIONS?(?: ADMINISTRATION HISTORY)?):?[\t \r]*\n
Medications Outside Hospital||(?:^[\t ]*MEDICATIONS? (?:AT )?OUTSIDE HOSPITAL):?[\t \r]*\n
Reason for Consult||(?:^[\t ]*REASON (?:FOR )?(?:CONSULT(?:ATION)?|REFERRAL)(?: ?\/? ?QUESTIONS?)?):?[\t \r]*\n
Problem List||(?:^[\t ]*(?:SIGNIFICANT )?PROBLEMS?(?: LIST)?):?[\t \r]*\n
Living Situation||(?:^[\t ]*LIV(?:E|ING) SITUATION):?[\t \r]*\n
Cytologic Diagnosis||(?:^[\t ]*CYTOLOGIC (?:DIAGNOSIS|DX)):?[\t \r]*\n
Discharge Instructions||(?:^[\t ]*DISCHARGE INSTRUCTIONS?):?[\t \r]*\n
Body Surface Area||(?:^[\t ]*(?:(?:BODY SURFACE AREA)|BSA)):?[\t \r]*\n
Discharge Condition||(?:^[\t ]*(?:(?:DISCHARGE CONDITION)|(?:CONDITION (?:(?:AT|ON) )?DISCHARGE))):?[\t \r]*\n
Diagnosis at Death||(?:^[\t ]*(?:(?:DIAGNOSIS|DX|CAUSE) (?:AT |OF )?DEATH)|COD):?[\t \r]*\n
Adverse Reactions||(?:^[\t ]*(?:(?:HISTORY (?:OF )?)?(?:ALLERG(?:Y|IES)|ADVERSE REACTIONS?))|(?:ALLERG(?:Y|IC|IES)(?: DISORDER)?(?:(?:\/| AND )ADVERSE REACTIONS?)?(?: HISTORY)?)):?[\t \r]*\n
