Numbered List||(?:^[\t ]*[\d]{1,2}(?::|\.)[\t ]+(?:(?!^[ ]*[\d]{1,2}(?::|\.)[\t ]+)(?:[^\t\r\n]+\r?\n))+){2,}||(?:^[\t ]*[\d]{1,2}(?::|\.)[\t ]+(?:(?!^[\t ]*[\d]{1,2}(?::|\.)[\t ]+)(?:[^\t\r\n]+\r?\n))+)
Alpha Sentence List||(?:^[\t ]*[A-Z](?::|\.)+\)?[\t ]+(?:[^\t\n\.]+(?:\.|\n))+\r?\n){2,}||(?:^[\t ]*[A-Z](?::|\.)+\)?[\t ]+(?:[^\t\n\.]+(?:\.|\n))+\r?\n)
Name Value List||(?:^[^\t\r\n]{2,50}:[\t ]+(?:[^\t\r\n:]+\r?\n)+){3,}||(?:^[^\t\r\n]{2,50}:[\t ]+(?:[^\t\r\n:]+\r?\n)+)
Multi Column List||(?:^(?:[^\t\r\n :]+(?: [^\t\r\n :]+)*(?:\t+| {3,}))+(?:[^\t\r\n ]+(?: [^\t\r\n ]+)*)[\t ]*\r?\n){3,}||\r?\n
// Mixed Column List||(?:^(?:[^\t\r\n :]+(?: [^\t\r\n :]+)*(?:\t+| {3,}))+(?:[^\t\r\n ]+(?: [^\t\r\n ]+)*)[\t ]*\r?\n[\t ]*(?:[^\t\r\n ]+(?: [^\t\r\n ]+)*)[\t ]*\r?\n){3,}||[\r\n][\t ]*(?:[^\t\r\n ]+(?: [^\t\r\n ]+)*)[\t ]*\r?\n
// Header List||(?:^[^\t\r\n\.]+\.{3,}[^\t\r\n\.]+\r?\n){3,}||\r?\n
Dash List||(?:^[\t ]*-{1,3}[\t ]+(?:(?:[^\t\r\n-]+-?)+\r?\n)+){2,}||(?:^[\t ]*-{1,3}[\t ]+(?:(?:[^\t\r\n-]+-?)+\r?\n)+)
Checkbox List||(?:^[\t ]*\[ *X? *\][^\r\n]+\r?\n){2,}||\r?\n
