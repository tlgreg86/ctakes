Identifying Data||(?:^[\t ]*IDENTIFYING DATA):?[\t \r]*\n
Chief Complaint||(?:^[\t ]*CHIEF COMPLAINT):?[\t \r]*\n
Clinical History||(?:^[\t ]*CLINICAL HISTORY):?[\t \r]*\n
Family History||(?:^[\t ]*FAMILY HISTORY):?[\t \r]*\n
History of Past Illness||(?:^[\t ]*(?:(?:HISTORY OF (?:THE )?PAST ILLNESS)|(?:PAST MEDICAL HISTORY))):?[\t \r]*\n
History of Present Illness||(?:^[\t ]*(?:HISTORY OF (?:THE )?(?:PRESENT|PHYSICAL) ILLNESS)(?: \(HPI(?:, PROBLEM BY PROBLEM)?\))?):?[\t \r]*\n
Current Health||(?:^[\t ]*CURRENT HEALTH(?: STATUS)?):?[\t \r]*\n
Psychosocial History||(?:^[\t ]*PSYCHOSOCIAL HISTORY):?[\t \r]*\n
Review of Systems||(?:^[\t ]*REVIEW OF SYSTEM)S?:?[\t \r]*\n
