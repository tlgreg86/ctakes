CUSTOM1|ctakes
CUSTOM1|ctakes application
CUSTOM2|new dictionary lookup
CUSTOM2|dictionary lookup, new
CUSTOM3|faster and stronger
CUSTOM3|stronger and faster

