CUSTOM1|APP1|ctakes
CUSTOM1|APP1|ctakes application
CUSTOM2|MOD1|new dictionary lookup
CUSTOM2|MOD1|dictionary lookup, new
CUSTOM3|DSC1|faster and stronger
CUSTOM3|DSC1|stronger and faster

