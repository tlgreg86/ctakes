1|19|claudition
2|21|pelvic
3|21|abdominal
4|109|aspirin
5|109|ibuprofen
6|109|acetaminophen
7|59|therapy
8|19|hyperlipidemia
9|109|supplement|dietary supplement
10|33|resting metabolic rate
11|21|knee
12|33|pain
13|21|colon
14|19|cancer
15|19|colon cancer
16|59|colonoscopy
17|33|discomfort
18|109|drug|pharmaceutical substance
19|21|arm
20|21|upper arm
21|33|swelling
22|59|arthroscopy
23|59|x-ray
24|33|shark bite
25|21|leg
26|109|narcotic
27|33|lesion
28|21|broca
